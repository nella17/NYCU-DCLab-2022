`timescale 1ns / 1ps
module lab9 (
    input clk,
    input reset_n,
    input [3:0] usr_btn,
    output LCD_RS,
    output LCD_RW,
    output LCD_E,
    output [3:0] LCD_D
);
endmodule
