`timescale 1ns / 1ps
module md5 (
    input  clk,
    input  reset_n,
    input  in,
    output reg out
);
endmodule
