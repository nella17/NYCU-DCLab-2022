`timescale 1ns / 1ps
module lab9_tb ();
endmodule
