`timescale 1ns / 1ps
/////////////////////////////////////////////////////////
module lab5(
    input clk,
    input reset_n,
    input [3:0] usr_btn,
    output [3:0] usr_led,
    output LCD_RS,
    output LCD_RW,
    output LCD_E,
    output [3:0] LCD_D
);

    // turn off all the LEDs
    assign usr_led = 4'b0000;

    wire btn_level, btn_pressed;
    reg prev_btn_level;
    reg [127:0] row_A = "Press BTN3 to   "; // Initialize the text of the first row. 
    reg [127:0] row_B = "show a message.."; // Initialize the text of the second row.

    LCD_module lcd0(
        .clk(clk),
        .reset(~reset_n),
        .row_A(row_A),
        .row_B(row_B),
        .LCD_E(LCD_E),
        .LCD_RS(LCD_RS),
        .LCD_RW(LCD_RW),
        .LCD_D(LCD_D)
    );

    debounce btn_db0(
        .clk(clk),
        .btn_input(usr_btn[3]),
        .btn_output(btn_level)
    );

    always @(posedge clk) begin
        if (~reset_n)
            prev_btn_level <= 1;
        else
            prev_btn_level <= btn_level;
    end

    assign btn_pressed = (btn_level == 1 && prev_btn_level == 0);

    always @(posedge clk) begin
        if (~reset_n) begin
            // Initialize the text when the user hit the reset button
            row_A = "Press BTN3 to   ";
            row_B = "show a message..";
        end else if (btn_pressed) begin
            row_A <= "Hello, World!   ";
            row_B <= "Demo of the LCD.";
        end
    end

endmodule

module debounce(
    input  clk,
    input  reset_n,
    input  in,
    output reg out
);
    reg init, stat;
    integer cnt;
    always @(posedge clk) begin
        if (!reset_n) begin
            init <= 0;
        end
        else begin
            if (init == 0 || stat != in) begin
                init <= 1;
                stat <= in;
                cnt <= 0;
            end
            else if (stat != out) begin
                if (cnt >= 10) begin
                    out <= stat;
                end
                cnt <= cnt+1;
            end
        end
    end
endmodule
